----------------------------------------------------------------------------------
-- Copyright (c) 2022 Burak Künkçü
-- Term Project - TermProjectLibrary (Library)
-- Character set mirrored from:
-- https://github.com/thelonious/vga_generator/blob/master/vga_text/font_rom.vhd
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;



package TermProjectLibrary is
function draw_char(X : natural; Y : natural; char : character) return boolean;
function draw_string(scanX : natural; scanY : natural; posX : natural; posY : natural; s : string; center : boolean; size : natural) return boolean;
function getStringRom1(index : natural) return String;
function getStringRom10(index : natural) return String;                                                        
function getStringRom100(index : natural) return String;
end TermProjectLibrary;


package body TermProjectLibrary is
function draw_char(X : natural; Y : natural; char : character) return boolean is

          constant ADDR_WIDTH: integer:=11;

          constant DATA_WIDTH: integer:=8;

          type rom_type is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);

         -- ROM definition

         constant ROM: rom_type:=(   -- 2^11-by-8

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "00000000", -- 5

         "00000000", -- 6

         "00000000", -- 7

         "00000000", -- 8

         "00000000", -- 9

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x01 ?

         "00000000", -- 0

         "00000000", -- 1

         "01111110", -- 2  ******

         "10000001", -- 3 *      *

         "10100101", -- 4 * *  * *

         "10000001", -- 5 *      *

         "10000001", -- 6 *      *

         "10111101", -- 7 * **** *

         "10011001", -- 8 *  **  *

         "10000001", -- 9 *      *

         "10000001", -- a *      *

         "01111110", -- b  ******

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x02 ?

         "00000000", -- 0

         "00000000", -- 1

         "01111110", -- 2  ******

         "11111111", -- 3 ********

         "11011011", -- 4 ** ** **

         "11111111", -- 5 ********

         "11111111", -- 6 ********

         "11000011", -- 7 **    **

         "11100111", -- 8 ***  ***

         "11111111", -- 9 ********

         "11111111", -- a ********

         "01111110", -- b  ******

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x03 ?

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "01101100", -- 4  ** **

         "11111110", -- 5 *******

         "11111110", -- 6 *******

         "11111110", -- 7 *******

         "11111110", -- 8 *******

         "01111100", -- 9  *****

         "00111000", -- a   ***

         "00010000", -- b    *

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x04 ?

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00010000", -- 4    *

         "00111000", -- 5   ***

         "01111100", -- 6  *****

         "11111110", -- 7 *******

         "01111100", -- 8  *****

         "00111000", -- 9   ***

         "00010000", -- a    *

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x05 ?

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00011000", -- 3    **

         "00111100", -- 4   ****

         "00111100", -- 5   ****

         "11100111", -- 6 ***  ***

         "11100111", -- 7 ***  ***

         "11100111", -- 8 ***  ***

         "00011000", -- 9    **

         "00011000", -- a    **

         "00111100", -- b   ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x06 ?

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00011000", -- 3    **

         "00111100", -- 4   ****

         "01111110", -- 5  ******

         "11111111", -- 6 ********

         "11111111", -- 7 ********

         "01111110", -- 8  ******

         "00011000", -- 9    **

         "00011000", -- a    **

         "00111100", -- b   ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x07 •

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "00000000", -- 5

         "00011000", -- 6    **

         "00111100", -- 7   ****

         "00111100", -- 8   ****

         "00011000", -- 9    **

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x08 ?

         "11111111", -- 0 ********

         "11111111", -- 1 ********

         "11111111", -- 2 ********

         "11111111", -- 3 ********

         "11111111", -- 4 ********

         "11111111", -- 5 ********

         "11100111", -- 6 ***  ***

         "11000011", -- 7 **    **

         "11000011", -- 8 **    **

         "11100111", -- 9 ***  ***

         "11111111", -- a ********

         "11111111", -- b ********

         "11111111", -- c ********

         "11111111", -- d ********

         "11111111", -- e ********

         "11111111", -- f ********

         -- code x09 ?

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "00111100", -- 5   ****

         "01100110", -- 6  **  **

         "01000010", -- 7  *    *

         "01000010", -- 8  *    *

         "01100110", -- 9  **  **

         "00111100", -- a   ****

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x0a ?

         "11111111", -- 0 ********

         "11111111", -- 1 ********

         "11111111", -- 2 ********

         "11111111", -- 3 ********

         "11111111", -- 4 ********

         "11000011", -- 5 **    **

         "10011001", -- 6 *  **  *

         "10111101", -- 7 * **** *

         "10111101", -- 8 * **** *

         "10011001", -- 9 *  **  *

         "11000011", -- a **    **

         "11111111", -- b ********

         "11111111", -- c ********

         "11111111", -- d ********

         "11111111", -- e ********

         "11111111", -- f ********

         -- code x0b ?

         "00000000", -- 0

         "00000000", -- 1

         "00011110", -- 2    ****

         "00001110", -- 3     ***

         "00011010", -- 4    ** *

         "00110010", -- 5   **  *

         "01111000", -- 6  ****

         "11001100", -- 7 **  **

         "11001100", -- 8 **  **

         "11001100", -- 9 **  **

         "11001100", -- a **  **

         "01111000", -- b  ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x0c ?

         "00000000", -- 0

         "00000000", -- 1

         "00111100", -- 2   ****

         "01100110", -- 3  **  **

         "01100110", -- 4  **  **

         "01100110", -- 5  **  **

         "01100110", -- 6  **  **

         "00111100", -- 7   ****

         "00011000", -- 8    **

         "01111110", -- 9  ******

         "00011000", -- a    **

         "00011000", -- b    **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x0d ?

         "00000000", -- 0

         "00000000", -- 1

         "00111111", -- 2   ******

         "00110011", -- 3   **  **

         "00111111", -- 4   ******

         "00110000", -- 5   **

         "00110000", -- 6   **

         "00110000", -- 7   **

         "00110000", -- 8   **

         "01110000", -- 9  ***

         "11110000", -- a ****

         "11100000", -- b ***

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x0e ?

         "00000000", -- 0

         "00000000", -- 1

         "01111111", -- 2  *******

         "01100011", -- 3  **   **

         "01111111", -- 4  *******

         "01100011", -- 5  **   **

         "01100011", -- 6  **   **

         "01100011", -- 7  **   **

         "01100011", -- 8  **   **

         "01100111", -- 9  **  ***

         "11100111", -- a ***  ***

         "11100110", -- b ***  **

         "11000000", -- c **

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x0f ?

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00011000", -- 3    **

         "00011000", -- 4    **

         "11011011", -- 5 ** ** **

         "00111100", -- 6   ****

         "11100111", -- 7 ***  ***

         "00111100", -- 8   ****

         "11011011", -- 9 ** ** **

         "00011000", -- a    **

         "00011000", -- b    **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x10 ?

         "00000000", -- 0

         "10000000", -- 1 *

         "11000000", -- 2 **

         "11100000", -- 3 ***

         "11110000", -- 4 ****

         "11111000", -- 5 *****

         "11111110", -- 6 *******

         "11111000", -- 7 *****

         "11110000", -- 8 ****

         "11100000", -- 9 ***

         "11000000", -- a **

         "10000000", -- b *

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x11 ?

         "00000000", -- 0

         "00000010", -- 1       *

         "00000110", -- 2      **

         "00001110", -- 3     ***

         "00011110", -- 4    ****

         "00111110", -- 5   *****

         "11111110", -- 6 *******

         "00111110", -- 7   *****

         "00011110", -- 8    ****

         "00001110", -- 9     ***

         "00000110", -- a      **

         "00000010", -- b       *

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x12 ?

         "00000000", -- 0

         "00000000", -- 1

         "00011000", -- 2    **

         "00111100", -- 3   ****

         "01111110", -- 4  ******

         "00011000", -- 5    **

         "00011000", -- 6    **

         "00011000", -- 7    **

         "01111110", -- 8  ******

         "00111100", -- 9   ****

         "00011000", -- a    **

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x13 ?

         "00000000", -- 0

         "00000000", -- 1

         "01100110", -- 2  **  **

         "01100110", -- 3  **  **

         "01100110", -- 4  **  **

         "01100110", -- 5  **  **

         "01100110", -- 6  **  **

         "01100110", -- 7  **  **

         "01100110", -- 8  **  **

         "00000000", -- 9

         "01100110", -- a  **  **

         "01100110", -- b  **  **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x14 ¶

         "00000000", -- 0

         "00000000", -- 1

         "01111111", -- 2  *******

         "11011011", -- 3 ** ** **

         "11011011", -- 4 ** ** **

         "11011011", -- 5 ** ** **

         "01111011", -- 6  **** **

         "00011011", -- 7    ** **

         "00011011", -- 8    ** **

         "00011011", -- 9    ** **

         "00011011", -- a    ** **

         "00011011", -- b    ** **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x15 §

         "00000000", -- 0

         "01111100", -- 1  *****

         "11000110", -- 2 **   **

         "01100000", -- 3  **

         "00111000", -- 4   ***

         "01101100", -- 5  ** **

         "11000110", -- 6 **   **

         "11000110", -- 7 **   **

         "01101100", -- 8  ** **

         "00111000", -- 9   ***

         "00001100", -- a     **

         "11000110", -- b **   **

         "01111100", -- c  *****

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x16 ?

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "00000000", -- 5

         "00000000", -- 6

         "00000000", -- 7

         "11111110", -- 8 *******

         "11111110", -- 9 *******

         "11111110", -- a *******

         "11111110", -- b *******

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x17 ?

         "00000000", -- 0

         "00000000", -- 1

         "00011000", -- 2    **

         "00111100", -- 3   ****

         "01111110", -- 4  ******

         "00011000", -- 5    **

         "00011000", -- 6    **

         "00011000", -- 7    **

         "01111110", -- 8  ******

         "00111100", -- 9   ****

         "00011000", -- a    **

         "01111110", -- b  ******

         "00110000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x18 ?

         "00000000", -- 0

         "00000000", -- 1

         "00011000", -- 2    **

         "00111100", -- 3   ****

         "01111110", -- 4  ******

         "00011000", -- 5    **

         "00011000", -- 6    **

         "00011000", -- 7    **

         "00011000", -- 8    **

         "00011000", -- 9    **

         "00011000", -- a    **

         "00011000", -- b    **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x19 ?

         "00000000", -- 0

         "00000000", -- 1

         "00011000", -- 2    **

         "00011000", -- 3    **

         "00011000", -- 4    **

         "00011000", -- 5    **

         "00011000", -- 6    **

         "00011000", -- 7    **

         "00011000", -- 8    **

         "01111110", -- 9  ******

         "00111100", -- a   ****

         "00011000", -- b    **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x1a ?

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "00011000", -- 5    **

         "00001100", -- 6     **

         "11111110", -- 7 *******

         "00001100", -- 8     **

         "00011000", -- 9    **

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x1b ?

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "00110000", -- 5   **

         "01100000", -- 6  **

         "11111110", -- 7 *******

         "01100000", -- 8  **

         "00110000", -- 9   **

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x1c ?

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "00000000", -- 5

         "11000000", -- 6 **

         "11000000", -- 7 **

         "11000000", -- 8 **

         "11111110", -- 9 *******

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x1d ?

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "00100100", -- 5   *  *

         "01100110", -- 6  **  **

         "11111111", -- 7 ********

         "01100110", -- 8  **  **

         "00100100", -- 9   *  *

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x1e ?

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00010000", -- 4    *

         "00111000", -- 5   ***

         "00111000", -- 6   ***

         "01111100", -- 7  *****

         "01111100", -- 8  *****

         "11111110", -- 9 *******

         "11111110", -- a *******

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x1f ?

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "11111110", -- 4 *******

         "11111110", -- 5 *******

         "01111100", -- 6  *****

         "01111100", -- 7  *****

         "00111000", -- 8   ***

         "00111000", -- 9   ***

         "00010000", -- a    *

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x20 ' '

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "00000000", -- 5

         "00000000", -- 6

         "00000000", -- 7

         "00000000", -- 8

         "00000000", -- 9

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x21 !

         "00000000", -- 0

         "00000000", -- 1

         "00011000", -- 2    **

         "00111100", -- 3   ****

         "00111100", -- 4   ****

         "00111100", -- 5   ****

         "00011000", -- 6    **

         "00011000", -- 7    **

         "00011000", -- 8    **

         "00000000", -- 9

         "00011000", -- a    **

         "00011000", -- b    **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x22 "

         "00000000", -- 0

         "01100110", -- 1  **  **

         "01100110", -- 2  **  **

         "01100110", -- 3  **  **

         "00100100", -- 4   *  *

         "00000000", -- 5

         "00000000", -- 6

         "00000000", -- 7

         "00000000", -- 8

         "00000000", -- 9

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x23 #

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "01101100", -- 3  ** **

         "01101100", -- 4  ** **

         "11111110", -- 5 *******

         "01101100", -- 6  ** **

         "01101100", -- 7  ** **

         "01101100", -- 8  ** **

         "11111110", -- 9 *******

         "01101100", -- a  ** **

         "01101100", -- b  ** **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x24 $

         "00011000", -- 0     **

         "00011000", -- 1     **

         "01111100", -- 2   *****

         "11000110", -- 3  **   **

         "11000010", -- 4  **    *

         "11000000", -- 5  **

         "01111100", -- 6   *****

         "00000110", -- 7       **

         "00000110", -- 8       **

         "10000110", -- 9  *    **

         "11000110", -- a  **   **

         "01111100", -- b   *****

         "00011000", -- c     **

         "00011000", -- d     **

         "00000000", -- e

         "00000000", -- f

         -- code x25 %

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "11000010", -- 4 **    *

         "11000110", -- 5 **   **

         "00001100", -- 6     **

         "00011000", -- 7    **

         "00110000", -- 8   **

         "01100000", -- 9  **

         "11000110", -- a **   **

         "10000110", -- b *    **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x26 &

         "00000000", -- 0

         "00000000", -- 1

         "00111000", -- 2   ***

         "01101100", -- 3  ** **

         "01101100", -- 4  ** **

         "00111000", -- 5   ***

         "01110110", -- 6  *** **

         "11011100", -- 7 ** ***

         "11001100", -- 8 **  **

         "11001100", -- 9 **  **

         "11001100", -- a **  **

         "01110110", -- b  *** **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x27 '

         "00000000", -- 0

         "00110000", -- 1   **

         "00110000", -- 2   **

         "00110000", -- 3   **

         "01100000", -- 4  **

         "00000000", -- 5

         "00000000", -- 6

         "00000000", -- 7

         "00000000", -- 8

         "00000000", -- 9

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x28 (

         "00000000", -- 0

         "00000000", -- 1

         "00001100", -- 2     **

         "00011000", -- 3    **

         "00110000", -- 4   **

         "00110000", -- 5   **

         "00110000", -- 6   **

         "00110000", -- 7   **

         "00110000", -- 8   **

         "00110000", -- 9   **

         "00011000", -- a    **

         "00001100", -- b     **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x29 )

         "00000000", -- 0

         "00000000", -- 1

         "00110000", -- 2   **

         "00011000", -- 3    **

         "00001100", -- 4     **

         "00001100", -- 5     **

         "00001100", -- 6     **

         "00001100", -- 7     **

         "00001100", -- 8     **

         "00001100", -- 9     **

         "00011000", -- a    **

         "00110000", -- b   **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x2a *

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "01100110", -- 5  **  **

         "00111100", -- 6   ****

         "11111111", -- 7 ********

         "00111100", -- 8   ****

         "01100110", -- 9  **  **

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x2b +

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "00011000", -- 5    **

         "00011000", -- 6    **

         "01111110", -- 7  ******

         "00011000", -- 8    **

         "00011000", -- 9    **

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x2c ,

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "00000000", -- 5

         "00000000", -- 6

         "00000000", -- 7

         "00000000", -- 8

         "00011000", -- 9    **

         "00011000", -- a    **

         "00011000", -- b    **

         "00110000", -- c   **

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x2d -

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "00000000", -- 5

         "00000000", -- 6

         "01111110", -- 7  ******

         "00000000", -- 8

         "00000000", -- 9

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x2e  .

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "00000000", -- 5

         "00000000", -- 6

         "00000000", -- 7

         "00000000", -- 8

         "00000000", -- 9

         "00011000", -- a    **

         "00011000", -- b    **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x2f /

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000010", -- 4       *

         "00000110", -- 5      **

         "00001100", -- 6     **

         "00011000", -- 7    **

         "00110000", -- 8   **

         "01100000", -- 9  **

         "11000000", -- a **

         "10000000", -- b *

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x30

         "00000000", -- 0

         "00000000", -- 1

         "01111100", -- 2  *****

         "11000110", -- 3 **   **

         "11000110", -- 4 **   **

         "11001110", -- 5 **  ***

         "11011110", -- 6 ** ****

         "11110110", -- 7 **** **

         "11100110", -- 8 ***  **

         "11000110", -- 9 **   **

         "11000110", -- a **   **

         "01111100", -- b  *****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x31 

         "00000000", -- 0

         "00000000", -- 1

         "00011000", -- 2

         "00111000", -- 3

         "01111000", -- 4    **

         "00011000", -- 5   ***

         "00011000", -- 6  ****

         "00011000", -- 7    **

         "00011000", -- 8    **

         "00011000", -- 9    **

         "00011000", -- a    **

         "01111110", -- b    **

         "00000000", -- c    **

         "00000000", -- d  ******

         "00000000", -- e

         "00000000", -- f

         -- code x32

         "00000000", -- 0

         "00000000", -- 1

         "01111100", -- 2  *****

         "11000110", -- 3 **   **

         "00000110", -- 4      **

         "00001100", -- 5     **

         "00011000", -- 6    **

         "00110000", -- 7   **

         "01100000", -- 8  **

         "11000000", -- 9 **

         "11000110", -- a **   **

         "11111110", -- b *******

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x33

         "00000000", -- 0

         "00000000", -- 1

         "01111100", -- 2  *****

         "11000110", -- 3 **   **

         "00000110", -- 4      **

         "00000110", -- 5      **

         "00111100", -- 6   ****

         "00000110", -- 7      **

         "00000110", -- 8      **

         "00000110", -- 9      **

         "11000110", -- a **   **

         "01111100", -- b  *****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x34

         "00000000", -- 0

         "00000000", -- 1

         "00001100", -- 2     **

         "00011100", -- 3    ***

         "00111100", -- 4   ****

         "01101100", -- 5  ** **

         "11001100", -- 6 **  **

         "11111110", -- 7 *******

         "00001100", -- 8     **

         "00001100", -- 9     **

         "00001100", -- a     **

         "00011110", -- b    ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x35

         "00000000", -- 0

         "00000000", -- 1

         "11111110", -- 2 *******

         "11000000", -- 3 **

         "11000000", -- 4 **

         "11000000", -- 5 **

         "11111100", -- 6 ******

         "00000110", -- 7      **

         "00000110", -- 8      **

         "00000110", -- 9      **

         "11000110", -- a **   **

         "01111100", -- b  *****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x36

         "00000000", -- 0

         "00000000", -- 1

         "00111000", -- 2   ***

         "01100000", -- 3  **

         "11000000", -- 4 **

         "11000000", -- 5 **

         "11111100", -- 6 ******

         "11000110", -- 7 **   **

         "11000110", -- 8 **   **

         "11000110", -- 9 **   **

         "11000110", -- a **   **

         "01111100", -- b  *****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x37

         "00000000", -- 0

         "00000000", -- 1

         "11111110", -- 2 *******

         "11000110", -- 3 **   **

         "00000110", -- 4      **

         "00000110", -- 5      **

         "00001100", -- 6     **

         "00011000", -- 7    **

         "00110000", -- 8   **

         "00110000", -- 9   **

         "00110000", -- a   **

         "00110000", -- b   **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x38

         "00000000", -- 0

         "00000000", -- 1

         "01111100", -- 2  *****

         "11000110", -- 3 **   **

         "11000110", -- 4 **   **

         "11000110", -- 5 **   **

         "01111100", -- 6  *****

         "11000110", -- 7 **   **

         "11000110", -- 8 **   **

         "11000110", -- 9 **   **

         "11000110", -- a **   **

         "01111100", -- b  *****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x39

         "00000000", -- 0

         "00000000", -- 1

         "01111100", -- 2  *****

         "11000110", -- 3 **   **

         "11000110", -- 4 **   **

         "11000110", -- 5 **   **

         "01111110", -- 6  ******

         "00000110", -- 7      **

         "00000110", -- 8      **

         "00000110", -- 9      **

         "00001100", -- a     **

         "01111000", -- b  ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x3a :

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00011000", -- 4    **

         "00011000", -- 5    **

         "00000000", -- 6

         "00000000", -- 7

         "00000000", -- 8

         "00011000", -- 9    **

         "00011000", -- a    **

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x3b ;

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00011000", -- 4    **

         "00011000", -- 5    **

         "00000000", -- 6

         "00000000", -- 7

         "00000000", -- 8

         "00011000", -- 9    **

         "00011000", -- a    **

         "00110000", -- b   **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x3c <

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000110", -- 3      **

         "00001100", -- 4     **

         "00011000", -- 5    **

         "00110000", -- 6   **

         "01100000", -- 7  **

         "00110000", -- 8   **

         "00011000", -- 9    **

         "00001100", -- a     **

         "00000110", -- b      **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x3d =

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "01111110", -- 5  ******

         "00000000", -- 6

         "00000000", -- 7

         "01111110", -- 8  ******

         "00000000", -- 9

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x3e >

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "01100000", -- 3  **

         "00110000", -- 4   **

         "00011000", -- 5    **

         "00001100", -- 6     **

         "00000110", -- 7      **

         "00001100", -- 8     **

         "00011000", -- 9    **

         "00110000", -- a   **

         "01100000", -- b  **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x3f ?

         "00000000", -- 0

         "00000000", -- 1

         "01111100", -- 2  *****

         "11000110", -- 3 **   **

         "11000110", -- 4 **   **

         "00001100", -- 5     **

         "00011000", -- 6    **

         "00011000", -- 7    **

         "00011000", -- 8    **

         "00000000", -- 9

         "00011000", -- a    **

         "00011000", -- b    **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x40 @

         "00000000", -- 0

         "00000000", -- 1

         "01111100", -- 2  *****

         "11000110", -- 3 **   **

         "11000110", -- 4 **   **

         "11000110", -- 5 **   **

         "11011110", -- 6 ** ****

         "11011110", -- 7 ** ****

         "11011110", -- 8 ** ****

         "11011100", -- 9 ** ***

         "11000000", -- a **

         "01111100", -- b  *****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x41

         "00000000", -- 0

         "00000000", -- 1

         "00010000", -- 2    *

         "00111000", -- 3   ***

         "01101100", -- 4  ** **

         "11000110", -- 5 **   **

         "11000110", -- 6 **   **

         "11111110", -- 7 *******

         "11000110", -- 8 **   **

         "11000110", -- 9 **   **

         "11000110", -- a **   **

         "11000110", -- b **   **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x42

         "00000000", -- 0

         "00000000", -- 1

         "11111100", -- 2 ******

         "01100110", -- 3  **  **

         "01100110", -- 4  **  **

         "01100110", -- 5  **  **

         "01111100", -- 6  *****

         "01100110", -- 7  **  **

         "01100110", -- 8  **  **

         "01100110", -- 9  **  **

         "01100110", -- a  **  **

         "11111100", -- b ******

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x43

         "00000000", -- 0

         "00000000", -- 1

         "00111100", -- 2   ****

         "01100110", -- 3  **  **

         "11000010", -- 4 **    *

         "11000000", -- 5 **

         "11000000", -- 6 **

         "11000000", -- 7 **

         "11000000", -- 8 **

         "11000010", -- 9 **    *

         "01100110", -- a  **  **

         "00111100", -- b   ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x44

         "00000000", -- 0

         "00000000", -- 1

         "11111000", -- 2 *****

         "01101100", -- 3  ** **

         "01100110", -- 4  **  **

         "01100110", -- 5  **  **

         "01100110", -- 6  **  **

         "01100110", -- 7  **  **

         "01100110", -- 8  **  **

         "01100110", -- 9  **  **

         "01101100", -- a  ** **

         "11111000", -- b *****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x45

         "00000000", -- 0

         "00000000", -- 1

         "11111110", -- 2 *******

         "01100110", -- 3  **  **

         "01100010", -- 4  **   *

         "01101000", -- 5  ** *

         "01111000", -- 6  ****

         "01101000", -- 7  ** *

         "01100000", -- 8  **

         "01100010", -- 9  **   *

         "01100110", -- a  **  **

         "11111110", -- b *******

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x46

         "00000000", -- 0

         "00000000", -- 1

         "11111110", -- 2 *******

         "01100110", -- 3  **  **

         "01100010", -- 4  **   *

         "01101000", -- 5  ** *

         "01111000", -- 6  ****

         "01101000", -- 7  ** *

         "01100000", -- 8  **

         "01100000", -- 9  **

         "01100000", -- a  **

         "11110000", -- b ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x47

         "00000000", -- 0

         "00000000", -- 1

         "00111100", -- 2   ****

         "01100110", -- 3  **  **

         "11000010", -- 4 **    *

         "11000000", -- 5 **

         "11000000", -- 6 **

         "11011110", -- 7 ** ****

         "11000110", -- 8 **   **

         "11000110", -- 9 **   **

         "01100110", -- a  **  **

         "00111010", -- b   *** *

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x48

         "00000000", -- 0

         "00000000", -- 1

         "11000110", -- 2 **   **

         "11000110", -- 3 **   **

         "11000110", -- 4 **   **

         "11000110", -- 5 **   **

         "11111110", -- 6 *******

         "11000110", -- 7 **   **

         "11000110", -- 8 **   **

         "11000110", -- 9 **   **

         "11000110", -- a **   **

         "11000110", -- b **   **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x49

         "00000000", -- 0

         "00000000", -- 1

         "00111100", -- 2   ****

         "00011000", -- 3    **

         "00011000", -- 4    **

         "00011000", -- 5    **

         "00011000", -- 6    **

         "00011000", -- 7    **

         "00011000", -- 8    **

         "00011000", -- 9    **

         "00011000", -- a    **

         "00111100", -- b   ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x4a

         "00000000", -- 0

         "00000000", -- 1

         "00011110", -- 2    ****

         "00001100", -- 3     **

         "00001100", -- 4     **

         "00001100", -- 5     **

         "00001100", -- 6     **

         "00001100", -- 7     **

         "11001100", -- 8 **  **

         "11001100", -- 9 **  **

         "11001100", -- a **  **

         "01111000", -- b  ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x4b

         "00000000", -- 0

         "00000000", -- 1

         "11100110", -- 2 ***  **

         "01100110", -- 3  **  **

         "01100110", -- 4  **  **

         "01101100", -- 5  ** **

         "01111000", -- 6  ****

         "01111000", -- 7  ****

         "01101100", -- 8  ** **

         "01100110", -- 9  **  **

         "01100110", -- a  **  **

         "11100110", -- b ***  **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x4c

         "00000000", -- 0

         "00000000", -- 1

         "11110000", -- 2 ****

         "01100000", -- 3  **

         "01100000", -- 4  **

         "01100000", -- 5  **

         "01100000", -- 6  **

         "01100000", -- 7  **

         "01100000", -- 8  **

         "01100010", -- 9  **   *

         "01100110", -- a  **  **

         "11111110", -- b *******

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x4d

         "00000000", -- 0

         "00000000", -- 1

         "11000011", -- 2 **    **

         "11100111", -- 3 ***  ***

         "11111111", -- 4 ********

         "11111111", -- 5 ********

         "11011011", -- 6 ** ** **

         "11000011", -- 7 **    **

         "11000011", -- 8 **    **

         "11000011", -- 9 **    **

         "11000011", -- a **    **

         "11000011", -- b **    **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x4e

         "00000000", -- 0

         "00000000", -- 1

         "11000110", -- 2 **   **

         "11100110", -- 3 ***  **

         "11110110", -- 4 **** **

         "11111110", -- 5 *******

         "11011110", -- 6 ** ****

         "11001110", -- 7 **  ***

         "11000110", -- 8 **   **

         "11000110", -- 9 **   **

         "11000110", -- a **   **

         "11000110", -- b **   **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x4f

         "00000000", -- 0

         "00000000", -- 1

         "01111100", -- 2  *****

         "11000110", -- 3 **   **

         "11000110", -- 4 **   **

         "11000110", -- 5 **   **

         "11000110", -- 6 **   **

         "11000110", -- 7 **   **

         "11000110", -- 8 **   **

         "11000110", -- 9 **   **

         "11000110", -- a **   **

         "01111100", -- b  *****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x50

         "00000000", -- 0

         "00000000", -- 1

         "11111100", -- 2 ******

         "01100110", -- 3  **  **

         "01100110", -- 4  **  **

         "01100110", -- 5  **  **

         "01111100", -- 6  *****

         "01100000", -- 7  **

         "01100000", -- 8  **

         "01100000", -- 9  **

         "01100000", -- a  **

         "11110000", -- b ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x510

         "00000000", -- 0

         "00000000", -- 1

         "01111100", -- 2  *****

         "11000110", -- 3 **   **

         "11000110", -- 4 **   **

         "11000110", -- 5 **   **

         "11000110", -- 6 **   **

         "11000110", -- 7 **   **

         "11000110", -- 8 **   **

         "11010110", -- 9 ** * **

         "11011110", -- a ** ****

         "01111100", -- b  *****

         "00001100", -- c     **

         "00001110", -- d     ***

         "00000000", -- e

         "00000000", -- f

         -- code x52

         "00000000", -- 0

         "00000000", -- 1

         "11111100", -- 2 ******

         "01100110", -- 3  **  **

         "01100110", -- 4  **  **

         "01100110", -- 5  **  **

         "01111100", -- 6  *****

         "01101100", -- 7  ** **

         "01100110", -- 8  **  **

         "01100110", -- 9  **  **

         "01100110", -- a  **  **

         "11100110", -- b ***  **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x53

         "00000000", -- 0

         "00000000", -- 1

         "01111100", -- 2  *****

         "11000110", -- 3 **   **

         "11000110", -- 4 **   **

         "01100000", -- 5  **

         "00111000", -- 6   ***

         "00001100", -- 7     **

         "00000110", -- 8      **

         "11000110", -- 9 **   **

         "11000110", -- a **   **

         "01111100", -- b  *****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x54

         "00000000", -- 0

         "00000000", -- 1

         "11111111", -- 2 ********

         "11011011", -- 3 ** ** **

         "10011001", -- 4 *  **  *

         "00011000", -- 5    **

         "00011000", -- 6    **

         "00011000", -- 7    **

         "00011000", -- 8    **

         "00011000", -- 9    **

         "00011000", -- a    **

         "00111100", -- b   ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x55

         "00000000", -- 0

         "00000000", -- 1

         "11000110", -- 2 **   **

         "11000110", -- 3 **   **

         "11000110", -- 4 **   **

         "11000110", -- 5 **   **

         "11000110", -- 6 **   **

         "11000110", -- 7 **   **

         "11000110", -- 8 **   **

         "11000110", -- 9 **   **

         "11000110", -- a **   **

         "01111100", -- b  *****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x56

         "00000000", -- 0

         "00000000", -- 1

         "11000011", -- 2 **    **

         "11000011", -- 3 **    **

         "11000011", -- 4 **    **

         "11000011", -- 5 **    **

         "11000011", -- 6 **    **

         "11000011", -- 7 **    **

         "11000011", -- 8 **    **

         "01100110", -- 9  **  **

         "00111100", -- a   ****

         "00011000", -- b    **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x57

         "00000000", -- 0

         "00000000", -- 1

         "11000011", -- 2 **    **

         "11000011", -- 3 **    **

         "11000011", -- 4 **    **

         "11000011", -- 5 **    **

         "11000011", -- 6 **    **

         "11011011", -- 7 ** ** **

         "11011011", -- 8 ** ** **

         "11111111", -- 9 ********

         "01100110", -- a  **  **

         "01100110", -- b  **  **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

      

         -- code x58

         "00000000", -- 0

         "00000000", -- 1

         "11000011", -- 2 **    **

         "11000011", -- 3 **    **

         "01100110", -- 4  **  **

         "00111100", -- 5   ****

         "00011000", -- 6    **

         "00011000", -- 7    **

         "00111100", -- 8   ****

         "01100110", -- 9  **  **

         "11000011", -- a **    **

         "11000011", -- b **    **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x59

         "00000000", -- 0

         "00000000", -- 1

         "11000011", -- 2 **    **

         "11000011", -- 3 **    **

         "11000011", -- 4 **    **

         "01100110", -- 5  **  **

         "00111100", -- 6   ****

         "00011000", -- 7    **

         "00011000", -- 8    **

         "00011000", -- 9    **

         "00011000", -- a    **

         "00111100", -- b   ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x5a

         "00000000", -- 0

         "00000000", -- 1

         "11111111", -- 2 ********

         "11000011", -- 3 **    **

         "10000110", -- 4 *    **

         "00001100", -- 5     **

         "00011000", -- 6    **

         "00110000", -- 7   **

         "01100000", -- 8  **

         "11000001", -- 9 **     *

         "11000011", -- a **    **

         "11111111", -- b ********

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x5b

         "00000000", -- 0

         "00000000", -- 1

         "00111100", -- 2   ****

         "00110000", -- 3   **

         "00110000", -- 4   **

         "00110000", -- 5   **

         "00110000", -- 6   **

         "00110000", -- 7   **

         "00110000", -- 8   **

         "00110000", -- 9   **

         "00110000", -- a   **

         "00111100", -- b   ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x5c

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "10000000", -- 3 *

         "11000000", -- 4 **

         "11100000", -- 5 ***

         "01110000", -- 6  ***

         "00111000", -- 7   ***

         "00011100", -- 8    ***

         "00001110", -- 9     ***

         "00000110", -- a      **

         "00000010", -- b       *

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x5d

         "00000000", -- 0

         "00000000", -- 1

         "00111100", -- 2   ****

         "00001100", -- 3     **

         "00001100", -- 4     **

         "00001100", -- 5     **

         "00001100", -- 6     **

         "00001100", -- 7     **

         "00001100", -- 8     **

         "00001100", -- 9     **

         "00001100", -- a     **

         "00111100", -- b   ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x5e

         "00010000", -- 0    *

         "00111000", -- 1   ***

         "01101100", -- 2  ** **

         "11000110", -- 3 **   **

         "00000000", -- 4

         "00000000", -- 5

         "00000000", -- 6

         "00000000", -- 7

         "00000000", -- 8

         "00000000", -- 9

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x5f

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "00000000", -- 5

         "00000000", -- 6

         "00000000", -- 7

         "00000000", -- 8

         "00000000", -- 9

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "11111111", -- d ********

         "00000000", -- e

         "00000000", -- f

         -- code x60

         "00110000", -- 0   **

         "00110000", -- 1   **

         "00011000", -- 2    **

         "00000000", -- 3

         "00000000", -- 4

         "00000000", -- 5

         "00000000", -- 6

         "00000000", -- 7

         "00000000", -- 8

         "00000000", -- 9

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x61

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "01111000", -- 5  ****

         "00001100", -- 6     **

         "01111100", -- 7  *****

         "11001100", -- 8 **  **

         "11001100", -- 9 **  **

         "11001100", -- a **  **

         "01110110", -- b  *** **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x62

         "00000000", -- 0

         "00000000", -- 1

         "11100000", -- 2  ***

         "01100000", -- 3   **

         "01100000", -- 4   **

         "01111000", -- 5   ****

         "01101100", -- 6   ** **

         "01100110", -- 7   **  **

         "01100110", -- 8   **  **

         "01100110", -- 9   **  **

         "01100110", -- a   **  **

         "01111100", -- b   *****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x63

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "01111100", -- 5  *****

         "11000110", -- 6 **   **

         "11000000", -- 7 **

         "11000000", -- 8 **

         "11000000", -- 9 **

         "11000110", -- a **   **

         "01111100", -- b  *****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x64

         "00000000", -- 0

         "00000000", -- 1

         "00011100", -- 2    ***

         "00001100", -- 3     **

         "00001100", -- 4     **

         "00111100", -- 5   ****

         "01101100", -- 6  ** **

         "11001100", -- 7 **  **

         "11001100", -- 8 **  **

         "11001100", -- 9 **  **

         "11001100", -- a **  **

         "01110110", -- b  *** **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x65

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "01111100", -- 5  *****

         "11000110", -- 6 **   **

         "11111110", -- 7 *******

         "11000000", -- 8 **

         "11000000", -- 9 **

         "11000110", -- a **   **

         "01111100", -- b  *****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x66

         "00000000", -- 0

         "00000000", -- 1

         "00111000", -- 2   ***

         "01101100", -- 3  ** **

         "01100100", -- 4  **  *

         "01100000", -- 5  **

         "11110000", -- 6 ****

         "01100000", -- 7  **

         "01100000", -- 8  **

         "01100000", -- 9  **

         "01100000", -- a  **

         "11110000", -- b ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x67

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "01110110", -- 5  *** **

         "11001100", -- 6 **  **

         "11001100", -- 7 **  **

         "11001100", -- 8 **  **

         "11001100", -- 9 **  **

         "11001100", -- a **  **

         "01111100", -- b  *****

         "00001100", -- c     **

         "11001100", -- d **  **

         "01111000", -- e  ****

         "00000000", -- f

         -- code x68

         "00000000", -- 0

         "00000000", -- 1

         "11100000", -- 2 ***

         "01100000", -- 3  **

         "01100000", -- 4  **

         "01101100", -- 5  ** **

         "01110110", -- 6  *** **

         "01100110", -- 7  **  **

         "01100110", -- 8  **  **

         "01100110", -- 9  **  **

         "01100110", -- a  **  **

         "11100110", -- b ***  **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x69

         "00000000", -- 0

         "00000000", -- 1

         "00011000", -- 2    **

         "00011000", -- 3    **

         "00000000", -- 4

         "00111000", -- 5   ***

         "00011000", -- 6    **

         "00011000", -- 7    **

         "00011000", -- 8    **

         "00011000", -- 9    **

         "00011000", -- a    **

         "00111100", -- b   ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x6a

         "00000000", -- 0

         "00000000", -- 1

         "00000110", -- 2      **

         "00000110", -- 3      **

         "00000000", -- 4

         "00001110", -- 5     ***

         "00000110", -- 6      **

         "00000110", -- 7      **

         "00000110", -- 8      **

         "00000110", -- 9      **

         "00000110", -- a      **

         "00000110", -- b      **

         "01100110", -- c  **  **

         "01100110", -- d  **  **

         "00111100", -- e   ****

         "00000000", -- f

         -- code x6b

         "00000000", -- 0

         "00000000", -- 1

         "11100000", -- 2 ***

         "01100000", -- 3  **

         "01100000", -- 4  **

         "01100110", -- 5  **  **

         "01101100", -- 6  ** **

         "01111000", -- 7  ****

         "01111000", -- 8  ****

         "01101100", -- 9  ** **

         "01100110", -- a  **  **

         "11100110", -- b ***  **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x6c

         "00000000", -- 0

         "00000000", -- 1

         "00111000", -- 2   ***

         "00011000", -- 3    **

         "00011000", -- 4    **

         "00011000", -- 5    **

         "00011000", -- 6    **

         "00011000", -- 7    **

         "00011000", -- 8    **

         "00011000", -- 9    **

         "00011000", -- a    **

         "00111100", -- b   ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x6d

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "11100110", -- 5 ***  **

         "11111111", -- 6 ********

         "11011011", -- 7 ** ** **

         "11011011", -- 8 ** ** **

         "11011011", -- 9 ** ** **

         "11011011", -- a ** ** **

         "11011011", -- b ** ** **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x6e

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "11011100", -- 5 ** ***

         "01100110", -- 6  **  **

         "01100110", -- 7  **  **

         "01100110", -- 8  **  **

         "01100110", -- 9  **  **

         "01100110", -- a  **  **

         "01100110", -- b  **  **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x6f

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "01111100", -- 5  *****

         "11000110", -- 6 **   **

         "11000110", -- 7 **   **

         "11000110", -- 8 **   **

         "11000110", -- 9 **   **

         "11000110", -- a **   **

         "01111100", -- b  *****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x70

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "11011100", -- 5 ** ***

         "01100110", -- 6  **  **

         "01100110", -- 7  **  **

         "01100110", -- 8  **  **

         "01100110", -- 9  **  **

         "01100110", -- a  **  **

         "01111100", -- b  *****

         "01100000", -- c  **

         "01100000", -- d  **

         "11110000", -- e ****

         "00000000", -- f

         -- code x71

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "01110110", -- 5  *** **

         "11001100", -- 6 **  **

         "11001100", -- 7 **  **

         "11001100", -- 8 **  **

         "11001100", -- 9 **  **

         "11001100", -- a **  **

         "01111100", -- b  *****

         "00001100", -- c     **

         "00001100", -- d     **

         "00011110", -- e    ****

         "00000000", -- f

         -- code x72

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "11011100", -- 5 ** ***

         "01110110", -- 6  *** **

         "01100110", -- 7  **  **

         "01100000", -- 8  **

         "01100000", -- 9  **

         "01100000", -- a  **

         "11110000", -- b ****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x73

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "01111100", -- 5  *****

         "11000110", -- 6 **   **

         "01100000", -- 7  **

         "00111000", -- 8   ***

         "00001100", -- 9     **

         "11000110", -- a **   **

         "01111100", -- b  *****

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x74

         "00000000", -- 0

         "00000000", -- 1

         "00010000", -- 2    *

         "00110000", -- 3   **

         "00110000", -- 4   **

         "11111100", -- 5 ******

         "00110000", -- 6   **

         "00110000", -- 7   **

         "00110000", -- 8   **

         "00110000", -- 9   **

         "00110110", -- a   ** **

         "00011100", -- b    ***

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x75

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "11001100", -- 5 **  **

         "11001100", -- 6 **  **

         "11001100", -- 7 **  **

         "11001100", -- 8 **  **

         "11001100", -- 9 **  **

         "11001100", -- a **  **

         "01110110", -- b  *** **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x76

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "11000011", -- 5 **    **

         "11000011", -- 6 **    **

         "11000011", -- 7 **    **

         "11000011", -- 8 **    **

         "01100110", -- 9  **  **

         "00111100", -- a   ****

         "00011000", -- b    **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x77

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "11000011", -- 5 **    **

         "11000011", -- 6 **    **

         "11000011", -- 7 **    **

         "11011011", -- 8 ** ** **

         "11011011", -- 9 ** ** **

         "11111111", -- a ********

         "01100110", -- b  **  **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x78

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "11000011", -- 5 **    **

         "01100110", -- 6  **  **

         "00111100", -- 7   ****

         "00011000", -- 8    **

         "00111100", -- 9   ****

         "01100110", -- a  **  **

         "11000011", -- b **    **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x79

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "11000110", -- 5 **   **

         "11000110", -- 6 **   **

         "11000110", -- 7 **   **

         "11000110", -- 8 **   **

         "11000110", -- 9 **   **

         "11000110", -- a **   **

         "01111110", -- b  ******

         "00000110", -- c      **

         "00001100", -- d     **

         "11111000", -- e *****

         "00000000", -- f

         -- code x7a

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00000000", -- 4

         "11111110", -- 5 *******

         "11001100", -- 6 **  **

         "00011000", -- 7    **

         "00110000", -- 8   **

         "01100000", -- 9  **

         "11000110", -- a **   **

         "11111110", -- b *******

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x7b {

         "00000000", -- 0

         "00000000", -- 1

         "00001110", -- 2     ***

         "00011000", -- 3    **

         "00011000", -- 4    **

         "00011000", -- 5    **

         "01110000", -- 6  ***

         "00011000", -- 7    **

         "00011000", -- 8    **

         "00011000", -- 9    **

         "00011000", -- a    **

         "00001110", -- b     ***

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x7c |

         "00000000", -- 0

         "00000000", -- 1

         "00011000", -- 2    **

         "00011000", -- 3    **

         "00011000", -- 4    **

         "00011000", -- 5    **

         "00000000", -- 6

         "00011000", -- 7    **

         "00011000", -- 8    **

         "00011000", -- 9    **

         "00011000", -- a    **

         "00011000", -- b    **

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x7d }

         "00000000", -- 0

         "00000000", -- 1

         "01110000", -- 2  ***

         "00011000", -- 3    **

         "00011000", -- 4    **

         "00011000", -- 5    **

         "00001110", -- 6     ***

         "00011000", -- 7    **

         "00011000", -- 8    **

         "00011000", -- 9    **

         "00011000", -- a    **

         "01110000", -- b  ***

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x7e ~

         "00000000", -- 0

         "00000000", -- 1

         "01110110", -- 2  *** **

         "11011100", -- 3 ** ***

         "00000000", -- 4

         "00000000", -- 5

         "00000000", -- 6

         "00000000", -- 7

         "00000000", -- 8

         "00000000", -- 9

         "00000000", -- a

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000", -- f

         -- code x7f

         "00000000", -- 0

         "00000000", -- 1

         "00000000", -- 2

         "00000000", -- 3

         "00010000", -- 4    *

         "00111000", -- 5   ***

         "01101100", -- 6  ** **

         "11000110", -- 7 **   **

         "11000110", -- 8 **   **

         "11000110", -- 9 **   **

         "11111110", -- a *******

         "00000000", -- b

         "00000000", -- c

         "00000000", -- d

         "00000000", -- e

         "00000000"  -- f

         );

      begin

          --return X <= 8 and Y <= 16 and ROM((char * 16) + Y)(9 - X) = '1';

          return ROM((CHARACTER'POS(char) * 16) + Y)(8 - X) = '1';

      end draw_char;

    

    function draw_string(scanX : natural; scanY : natural; posX : natural; posY : natural; s : string; center : boolean; size : natural) return boolean is

    constant charW : natural := 8 * size;

    constant charWsp : natural := charW + 2;

    constant charH : natural := 16 * size;

    constant width : natural := charWsp * s'LENGTH;

    constant height : natural := charH;

    variable x : natural := posX;

    variable y : natural := posY;

    variable char : natural;

    variable subX : natural;

    begin

        if (center) then

            x := x - (width / 2);

            y := y - (height / 2);

         end if;

  

         if (scanX < x or scanY < y) then

             return false;

         end if;

      

         if (scanX - x > width or scanY - y > height) then

             return false;

         end if;

      

         x := scanX - x;

         y := scanY - y;

      

         subX := x mod charWsp;

         char := (x / charWsp) + 1;

      

         return draw_char(subX / size, y / size, s(char));

    end draw_string;   

    

    function getStringRom1(index : natural) return String is

    type StringRomType1 is array(0 to 9) of String(1 to 1);

    constant StringRom1 : StringRomType1 := (0 => "0", 1 => "1", 2 => "2", 3 => "3", 4 => "4", 5 => "5", 6 => "6", 7 => "7", 8 => "8", 9 => "9");

    begin

        return StringRom1(index mod 10);

    end getStringRom1;

    

    function getStringRom10(index : natural) return String is

    type StringRomType10 is array(10 to 99) of String(1 to 2);

    constant StringRom10 : StringRomType10 := (10 => "10", 11 => "11", 12 => "12", 13 => "13", 14 => "14", 15 => "15", 16 => "16", 17 => "17", 

        18 => "18", 19 => "19", 20 => "20", 21 => "21", 22 => "22", 23 => "23", 24 => "24", 25 => "25", 26 => "26", 27 => "27", 28 => "28", 

        29 => "29", 30 => "30", 31 => "31", 32 => "32", 33 => "33", 34 => "34", 35 => "35", 36 => "36", 37 => "37", 38 => "38", 39 => "39",

        40 => "40", 41 => "41", 42 => "42", 43 => "43", 44 => "44", 45 => "45", 46 => "46", 47 => "47", 48 => "48", 49 => "49", 50 => "50", 

        51 => "51", 52 => "52", 53 => "53", 54 => "54", 55 => "55", 56 => "56", 57 => "57", 58 => "58", 59 => "59", 60 => "60", 61 => "61", 

        62 => "62", 63 => "63", 64 => "64", 65 => "65", 66 => "66", 67 => "67", 68 => "68", 69 => "69", 70 => "70", 71 => "71", 72 => "72", 

        73 => "73", 74 => "74", 75 => "75", 76 => "76", 77 => "77", 78 => "78", 79 => "79", 80 => "80", 81 => "81", 82 => "82", 83 => "83", 

        84 => "84", 85 => "85", 86 => "86", 87 => "87", 88 => "88", 89 => "89", 90 => "90", 91 => "91", 92 => "92", 93 => "93", 94 => "94", 

        95 => "95", 96 => "96", 97 => "97", 98 => "98", 99 => "99");

    begin

        return StringRom10(index mod 100);

    end getStringRom10;

    

    function getStringRom100(index : natural) return String is

    type StringRomType100 is array(100 to 999) of String(1 to 3);

    constant StringRom100 : StringRomType100 := (100 => "100", 101 => "101", 102 => "102", 103 => "103", 104 => "104", 105 => "105", 106 => "106",

        107 => "107", 108 => "108", 109 => "109", 110 => "110", 111 => "111", 112 => "112", 113 => "113", 114 => "114", 115 => "115", 116 => "116",

        117 => "117", 118 => "118", 119 => "119", 120 => "120", 121 => "121", 122 => "122", 123 => "123", 124 => "124", 125 => "125", 126 => "126",

        127 => "127", 128 => "128", 129 => "129", 130 => "130", 131 => "131", 132 => "132", 133 => "133", 134 => "134", 135 => "135", 136 => "136",

        137 => "137", 138 => "138", 139 => "139", 140 => "140", 141 => "141", 142 => "142", 143 => "143", 144 => "144", 145 => "145", 146 => "146", 

        147 => "147", 148 => "148", 149 => "149", 150 => "150", 151 => "151", 152 => "152", 153 => "153", 154 => "154", 155 => "155", 156 => "156", 

        157 => "157", 158 => "158", 159 => "159", 160 => "160", 161 => "161", 162 => "162", 163 => "163", 164 => "164", 165 => "165", 166 => "166", 

        167 => "167", 168 => "168", 169 => "169", 170 => "170", 171 => "171", 172 => "172", 173 => "173", 174 => "174", 175 => "175", 176 => "176", 

        177 => "177", 178 => "178", 179 => "179", 180 => "180", 181 => "181", 182 => "182", 183 => "183", 184 => "184", 185 => "185", 186 => "186", 

        187 => "187", 188 => "188", 189 => "189", 190 => "190", 191 => "191", 192 => "192", 193 => "193", 194 => "194", 195 => "195", 196 => "196", 

        197 => "197", 198 => "198", 199 => "199", 200 => "200", 201 => "201", 202 => "202", 203 => "203", 204 => "204", 205 => "205", 206 => "206", 

        207 => "207", 208 => "208", 209 => "209", 210 => "210", 211 => "211", 212 => "212", 213 => "213", 214 => "214", 215 => "215", 216 => "216",

        217 => "217", 218 => "218", 219 => "219", 220 => "220", 221 => "221", 222 => "222", 223 => "223", 224 => "224", 225 => "225", 226 => "226",

        227 => "227", 228 => "228", 229 => "229", 230 => "230", 231 => "231", 232 => "232", 233 => "233", 234 => "234", 235 => "235", 236 => "236", 

        237 => "237", 238 => "238", 239 => "239", 240 => "240", 241 => "241", 242 => "242", 243 => "243", 244 => "244", 245 => "245", 246 => "246",

        247 => "247", 248 => "248", 249 => "249", 250 => "250", 251 => "251", 252 => "252", 253 => "253", 254 => "254", 255 => "255", 256 => "256",

        257 => "257", 258 => "258", 259 => "259", 260 => "260", 261 => "261", 262 => "262", 263 => "263", 264 => "264", 265 => "265", 266 => "266",

        267 => "267", 268 => "268", 269 => "269", 270 => "270", 271 => "271", 272 => "272", 273 => "273", 274 => "274", 275 => "275", 276 => "276",

        277 => "277", 278 => "278", 279 => "279", 280 => "280", 281 => "281", 282 => "282", 283 => "283", 284 => "284", 285 => "285", 286 => "286", 

        287 => "287", 288 => "288", 289 => "289", 290 => "290", 291 => "291", 292 => "292", 293 => "293", 294 => "294", 295 => "295", 296 => "296", 

        297 => "297", 298 => "298", 299 => "299", 300 => "300", 301 => "301", 302 => "302", 303 => "303", 304 => "304", 305 => "305", 306 => "306",

        307 => "307", 308 => "308", 309 => "309", 310 => "310", 311 => "311", 312 => "312", 313 => "313", 314 => "314", 315 => "315", 316 => "316",

        317 => "317", 318 => "318", 319 => "319", 320 => "320", 321 => "321", 322 => "322", 323 => "323", 324 => "324", 325 => "325", 326 => "326", 

        327 => "327", 328 => "328", 329 => "329", 330 => "330", 331 => "331", 332 => "332", 333 => "333", 334 => "334", 335 => "335", 336 => "336",

        337 => "337", 338 => "338", 339 => "339", 340 => "340", 341 => "341", 342 => "342", 343 => "343", 344 => "344", 345 => "345", 346 => "346", 

        347 => "347", 348 => "348", 349 => "349", 350 => "350", 351 => "351", 352 => "352", 353 => "353", 354 => "354", 355 => "355", 356 => "356", 

        357 => "357", 358 => "358", 359 => "359", 360 => "360", 361 => "361", 362 => "362", 363 => "363", 364 => "364", 365 => "365", 366 => "366", 

        367 => "367", 368 => "368", 369 => "369", 370 => "370", 371 => "371", 372 => "372", 373 => "373", 374 => "374", 375 => "375", 376 => "376", 

        377 => "377", 378 => "378", 379 => "379", 380 => "380", 381 => "381", 382 => "382", 383 => "383", 384 => "384", 385 => "385", 386 => "386",

        387 => "387", 388 => "388", 389 => "389", 390 => "390", 391 => "391", 392 => "392", 393 => "393", 394 => "394", 395 => "395", 396 => "396",

        397 => "397", 398 => "398", 399 => "399", 400 => "400", 401 => "401", 402 => "402", 403 => "403", 404 => "404", 405 => "405", 406 => "406",

        407 => "407", 408 => "408", 409 => "409", 410 => "410", 411 => "411", 412 => "412", 413 => "413", 414 => "414", 415 => "415", 416 => "416", 

        417 => "417", 418 => "418", 419 => "419", 420 => "420", 421 => "421", 422 => "422", 423 => "423", 424 => "424", 425 => "425", 426 => "426", 

        427 => "427", 428 => "428", 429 => "429", 430 => "430", 431 => "431", 432 => "432", 433 => "433", 434 => "434", 435 => "435", 436 => "436", 

        437 => "437", 438 => "438", 439 => "439", 440 => "440", 441 => "441", 442 => "442", 443 => "443", 444 => "444", 445 => "445", 446 => "446", 

        447 => "447", 448 => "448", 449 => "449", 450 => "450", 451 => "451", 452 => "452", 453 => "453", 454 => "454", 455 => "455", 456 => "456", 

        457 => "457", 458 => "458", 459 => "459", 460 => "460", 461 => "461", 462 => "462", 463 => "463", 464 => "464", 465 => "465", 466 => "466", 

        467 => "467", 468 => "468", 469 => "469", 470 => "470", 471 => "471", 472 => "472", 473 => "473", 474 => "474", 475 => "475", 476 => "476", 

        477 => "477", 478 => "478", 479 => "479", 480 => "480", 481 => "481", 482 => "482", 483 => "483", 484 => "484", 485 => "485", 486 => "486", 

        487 => "487", 488 => "488", 489 => "489", 490 => "490", 491 => "491", 492 => "492", 493 => "493", 494 => "494", 495 => "495", 496 => "496", 

        497 => "497", 498 => "498", 499 => "499", 500 => "500", 501 => "501", 502 => "502", 503 => "503", 504 => "504", 505 => "505", 506 => "506", 

        507 => "507", 508 => "508", 509 => "509", 510 => "510", 511 => "511", 512 => "512", 513 => "513", 514 => "514", 515 => "515", 516 => "516", 

        517 => "517", 518 => "518", 519 => "519", 520 => "520", 521 => "521", 522 => "522", 523 => "523", 524 => "524", 525 => "525", 526 => "526", 

        527 => "527", 528 => "528", 529 => "529", 530 => "530", 531 => "531", 532 => "532", 533 => "533", 534 => "534", 535 => "535", 536 => "536", 

        537 => "537", 538 => "538", 539 => "539", 540 => "540", 541 => "541", 542 => "542", 543 => "543", 544 => "544", 545 => "545", 546 => "546", 

        547 => "547", 548 => "548", 549 => "549", 550 => "550", 551 => "551", 552 => "552", 553 => "553", 554 => "554", 555 => "555", 556 => "556", 

        557 => "557", 558 => "558", 559 => "559", 560 => "560", 561 => "561", 562 => "562", 563 => "563", 564 => "564", 565 => "565", 566 => "566", 

        567 => "567", 568 => "568", 569 => "569", 570 => "570", 571 => "571", 572 => "572", 573 => "573", 574 => "574", 575 => "575", 576 => "576", 

        577 => "577", 578 => "578", 579 => "579", 580 => "580", 581 => "581", 582 => "582", 583 => "583", 584 => "584", 585 => "585", 586 => "586", 

        587 => "587", 588 => "588", 589 => "589", 590 => "590", 591 => "591", 592 => "592", 593 => "593", 594 => "594", 595 => "595", 596 => "596", 

        597 => "597", 598 => "598", 599 => "599", 600 => "600", 601 => "601", 602 => "602", 603 => "603", 604 => "604", 605 => "605", 606 => "606", 

        607 => "607", 608 => "608", 609 => "609", 610 => "610", 611 => "611", 612 => "612", 613 => "613", 614 => "614", 615 => "615", 616 => "616", 

        617 => "617", 618 => "618", 619 => "619", 620 => "620", 621 => "621", 622 => "622", 623 => "623", 624 => "624", 625 => "625", 626 => "626", 

        627 => "627", 628 => "628", 629 => "629", 630 => "630", 631 => "631", 632 => "632", 633 => "633", 634 => "634", 635 => "635", 636 => "636", 

        637 => "637", 638 => "638", 639 => "639", 640 => "640", 641 => "641", 642 => "642", 643 => "643", 644 => "644", 645 => "645", 646 => "646", 

        647 => "647", 648 => "648", 649 => "649", 650 => "650", 651 => "651", 652 => "652", 653 => "653", 654 => "654", 655 => "655", 656 => "656", 

        657 => "657", 658 => "658", 659 => "659", 660 => "660", 661 => "661", 662 => "662", 663 => "663", 664 => "664", 665 => "665", 666 => "666", 

        667 => "667", 668 => "668", 669 => "669", 670 => "670", 671 => "671", 672 => "672", 673 => "673", 674 => "674", 675 => "675", 676 => "676", 

        677 => "677", 678 => "678", 679 => "679", 680 => "680", 681 => "681", 682 => "682", 683 => "683", 684 => "684", 685 => "685", 686 => "686", 

        687 => "687", 688 => "688", 689 => "689", 690 => "690", 691 => "691", 692 => "692", 693 => "693", 694 => "694", 695 => "695", 696 => "696", 

        697 => "697", 698 => "698", 699 => "699", 700 => "700", 701 => "701", 702 => "702", 703 => "703", 704 => "704", 705 => "705", 706 => "706", 

        707 => "707", 708 => "708", 709 => "709", 710 => "710", 711 => "711", 712 => "712", 713 => "713", 714 => "714", 715 => "715", 716 => "716", 

        717 => "717", 718 => "718", 719 => "719", 720 => "720", 721 => "721", 722 => "722", 723 => "723", 724 => "724", 725 => "725", 726 => "726", 

        727 => "727", 728 => "728", 729 => "729", 730 => "730", 731 => "731", 732 => "732", 733 => "733", 734 => "734", 735 => "735", 736 => "736", 

        737 => "737", 738 => "738", 739 => "739", 740 => "740", 741 => "741", 742 => "742", 743 => "743", 744 => "744", 745 => "745", 746 => "746", 

        747 => "747", 748 => "748", 749 => "749", 750 => "750", 751 => "751", 752 => "752", 753 => "753", 754 => "754", 755 => "755", 756 => "756", 

        757 => "757", 758 => "758", 759 => "759", 760 => "760", 761 => "761", 762 => "762", 763 => "763", 764 => "764", 765 => "765", 766 => "766", 

        767 => "767", 768 => "768", 769 => "769", 770 => "770", 771 => "771", 772 => "772", 773 => "773", 774 => "774", 775 => "775", 776 => "776", 

        777 => "777", 778 => "778", 779 => "779", 780 => "780", 781 => "781", 782 => "782", 783 => "783", 784 => "784", 785 => "785", 786 => "786", 

        787 => "787", 788 => "788", 789 => "789", 790 => "790", 791 => "791", 792 => "792", 793 => "793", 794 => "794", 795 => "795", 796 => "796", 

        797 => "797", 798 => "798", 799 => "799", 800 => "800", 801 => "801", 802 => "802", 803 => "803", 804 => "804", 805 => "805", 806 => "806", 

        807 => "807", 808 => "808", 809 => "809", 810 => "810", 811 => "811", 812 => "812", 813 => "813", 814 => "814", 815 => "815", 816 => "816", 

        817 => "817", 818 => "818", 819 => "819", 820 => "820", 821 => "821", 822 => "822", 823 => "823", 824 => "824", 825 => "825", 826 => "826", 

        827 => "827", 828 => "828", 829 => "829", 830 => "830", 831 => "831", 832 => "832", 833 => "833", 834 => "834", 835 => "835", 836 => "836", 

        837 => "837", 838 => "838", 839 => "839", 840 => "840", 841 => "841", 842 => "842", 843 => "843", 844 => "844", 845 => "845", 846 => "846", 

        847 => "847", 848 => "848", 849 => "849", 850 => "850", 851 => "851", 852 => "852", 853 => "853", 854 => "854", 855 => "855", 856 => "856", 

        857 => "857", 858 => "858", 859 => "859", 860 => "860", 861 => "861", 862 => "862", 863 => "863", 864 => "864", 865 => "865", 866 => "866", 

        867 => "867", 868 => "868", 869 => "869", 870 => "870", 871 => "871", 872 => "872", 873 => "873", 874 => "874", 875 => "875", 876 => "876", 

        877 => "877", 878 => "878", 879 => "879", 880 => "880", 881 => "881", 882 => "882", 883 => "883", 884 => "884", 885 => "885", 886 => "886", 

        887 => "887", 888 => "888", 889 => "889", 890 => "890", 891 => "891", 892 => "892", 893 => "893", 894 => "894", 895 => "895", 896 => "896", 

        897 => "897", 898 => "898", 899 => "899", 900 => "900", 901 => "901", 902 => "902", 903 => "903", 904 => "904", 905 => "905", 906 => "906", 

        907 => "907", 908 => "908", 909 => "909", 910 => "910", 911 => "911", 912 => "912", 913 => "913", 914 => "914", 915 => "915", 916 => "916", 

        917 => "917", 918 => "918", 919 => "919", 920 => "920", 921 => "921", 922 => "922", 923 => "923", 924 => "924", 925 => "925", 926 => "926", 

        927 => "927", 928 => "928", 929 => "929", 930 => "930", 931 => "931", 932 => "932", 933 => "933", 934 => "934", 935 => "935", 936 => "936", 

        937 => "937", 938 => "938", 939 => "939", 940 => "940", 941 => "941", 942 => "942", 943 => "943", 944 => "944", 945 => "945", 946 => "946", 

        947 => "947", 948 => "948", 949 => "949", 950 => "950", 951 => "951", 952 => "952", 953 => "953", 954 => "954", 955 => "955", 956 => "956", 

        957 => "957", 958 => "958", 959 => "959", 960 => "960", 961 => "961", 962 => "962", 963 => "963", 964 => "964", 965 => "965", 966 => "966", 

        967 => "967", 968 => "968", 969 => "969", 970 => "970", 971 => "971", 972 => "972", 973 => "973", 974 => "974", 975 => "975", 976 => "976", 

        977 => "977", 978 => "978", 979 => "979", 980 => "980", 981 => "981", 982 => "982", 983 => "983", 984 => "984", 985 => "985", 986 => "986", 

        987 => "987", 988 => "988", 989 => "989", 990 => "990", 991 => "991", 992 => "992", 993 => "993", 994 => "994", 995 => "995", 996 => "996", 

        997 => "997", 998 => "998", 999 => "999");

    begin

        return StringRom100(index mod 1000);

    end getStringRom100;

end TermProjectLibrary;